netcdf LHM_ZW_LHM_MozartDistrict_REF2017BP18 {
dimensions:
	analysis_time = 1 ;
	stations = 244 ;
	string64 = 64 ;
	string255 = 255 ;
	time = 3636 ;
variables:
	double analysis_time(analysis_time) ;
		analysis_time:_FillValue = NaN ;
		analysis_time:standard_name = "forecast_reference_time" ;
		analysis_time:long_name = "forecast_reference_time" ;
		analysis_time:units = "minutes since 1970-01-01T00:00:00+00:00" ;
		analysis_time:calendar = "proleptic_gregorian" ;
	double lat(stations) ;
		lat:_FillValue = 9.96921e+36 ;
		lat:standard_name = "latitude" ;
		lat:long_name = "Station coordinates, latitude" ;
		lat:units = "degrees_north" ;
		lat:axis = "Y" ;
	double lon(stations) ;
		lon:_FillValue = 9.96921e+36 ;
		lon:standard_name = "longitude" ;
		lon:long_name = "Station coordinates, longitude" ;
		lon:units = "degrees_east" ;
		lon:axis = "X" ;
	double y(stations) ;
		y:_FillValue = 9.96921e+36 ;
		y:standard_name = "projection_y_coordinate" ;
		y:long_name = "y coordinate according to Rijks Driehoekstelsel" ;
		y:units = "m" ;
		y:axis = "Y" ;
		y:coordinates = "lon lat" ;
	double x(stations) ;
		x:_FillValue = 9.96921e+36 ;
		x:standard_name = "projection_x_coordinate" ;
		x:long_name = "x coordinate according to Rijks Driehoekstelsel" ;
		x:units = "m" ;
		x:axis = "X" ;
		x:coordinates = "lon lat" ;
	double z(stations) ;
		z:_FillValue = 9.96921e+36 ;
		z:long_name = "height above mean sea level" ;
		z:units = "meters" ;
		z:coordinates = "lon lat" ;
	char station_id(stations, string64) ;
		station_id:long_name = "station identification code" ;
		station_id:cf_role = "timeseries_id" ;
		station_id:coordinates = "lon lat" ;
	char station_names(stations, string255) ;
		station_names:long_name = "station name" ;
		station_names:coordinates = "lon lat" ;
	int64 time(time) ;
		time:standard_name = "time" ;
		time:long_name = "time" ;
		time:axis = "T" ;
		time:units = "days since 1911-01-11 00:00:00" ;
		time:calendar = "proleptic_gregorian" ;
	float precip(time, stations) ;
		precip:_FillValue = -999.f ;
		precip:long_name = "precip" ;
		precip:units = "m3" ;
		precip:coordinates = "lon lat" ;
	float evaporation(time, stations) ;
		evaporation:_FillValue = -999.f ;
		evaporation:long_name = "evaporation" ;
		evaporation:units = "m3" ;
		evaporation:coordinates = "lon lat" ;
	float drainage_sh(time, stations) ;
		drainage_sh:_FillValue = -999.f ;
		drainage_sh:long_name = "drainage_sh" ;
		drainage_sh:units = "m3" ;
		drainage_sh:coordinates = "lon lat" ;
	float drainage_dp(time, stations) ;
		drainage_dp:_FillValue = -999.f ;
		drainage_dp:long_name = "drainage_dp" ;
		drainage_dp:units = "m3" ;
		drainage_dp:coordinates = "lon lat" ;
	float infiltration_sh(time, stations) ;
		infiltration_sh:_FillValue = -999.f ;
		infiltration_sh:long_name = "infiltration_sh" ;
		infiltration_sh:units = "m3" ;
		infiltration_sh:coordinates = "lon lat" ;
	byte infiltration_dp(time, stations) ;
		infiltration_dp:_FillValue = -128b ;
		infiltration_dp:long_name = "infiltration_dp" ;
		infiltration_dp:units = "m3" ;
		infiltration_dp:coordinates = "lon lat" ;
		infiltration_dp:add_offset = 0.f ;
		infiltration_dp:scale_factor = 0.01f ;
	float urbanrunoff(time, stations) ;
		urbanrunoff:_FillValue = -999.f ;
		urbanrunoff:long_name = "urbanrunoff" ;
		urbanrunoff:units = "m3" ;
		urbanrunoff:coordinates = "lon lat" ;
	float upstream(time, stations) ;
		upstream:_FillValue = -999.f ;
		upstream:long_name = "upstream" ;
		upstream:units = "m3" ;
		upstream:coordinates = "lon lat" ;
	float downstream(time, stations) ;
		downstream:_FillValue = -999.f ;
		downstream:long_name = "downstream" ;
		downstream:units = "m3" ;
		downstream:coordinates = "lon lat" ;
	float from_dw(time, stations) ;
		from_dw:_FillValue = -999.f ;
		from_dw:long_name = "from_dw" ;
		from_dw:units = "m3" ;
		from_dw:coordinates = "lon lat" ;
	float to_dw(time, stations) ;
		to_dw:_FillValue = -999.f ;
		to_dw:long_name = "to_dw" ;
		to_dw:units = "m3" ;
		to_dw:coordinates = "lon lat" ;
	float dstorage(time, stations) ;
		dstorage:_FillValue = -999.f ;
		dstorage:long_name = "dstorage" ;
		dstorage:units = "m3" ;
		dstorage:coordinates = "lon lat" ;
	float alloc_agric(time, stations) ;
		alloc_agric:_FillValue = -999.f ;
		alloc_agric:long_name = "alloc_agric" ;
		alloc_agric:units = "m3" ;
		alloc_agric:coordinates = "lon lat" ;
	float alloc_wm(time, stations) ;
		alloc_wm:_FillValue = -999.f ;
		alloc_wm:long_name = "alloc_wm" ;
		alloc_wm:units = "m3" ;
		alloc_wm:coordinates = "lon lat" ;
	float alloc_flush(time, stations) ;
		alloc_flush:_FillValue = -999.f ;
		alloc_flush:long_name = "alloc_flush" ;
		alloc_flush:units = "m3" ;
		alloc_flush:coordinates = "lon lat" ;
	float alloc_flushreturn(time, stations) ;
		alloc_flushreturn:_FillValue = -999.f ;
		alloc_flushreturn:long_name = "alloc_flushreturn" ;
		alloc_flushreturn:units = "m3" ;
		alloc_flushreturn:coordinates = "lon lat" ;
	byte alloc_pubwat(time, stations) ;
		alloc_pubwat:_FillValue = -128b ;
		alloc_pubwat:long_name = "alloc_pubwat" ;
		alloc_pubwat:units = "m3" ;
		alloc_pubwat:coordinates = "lon lat" ;
		alloc_pubwat:add_offset = 0.f ;
		alloc_pubwat:scale_factor = 0.01f ;
	byte alloc_industry(time, stations) ;
		alloc_industry:_FillValue = -128b ;
		alloc_industry:long_name = "alloc_industry" ;
		alloc_industry:units = "m3" ;
		alloc_industry:coordinates = "lon lat" ;
		alloc_industry:add_offset = 0.f ;
		alloc_industry:scale_factor = 0.01f ;
	byte alloc_greenhouse(time, stations) ;
		alloc_greenhouse:_FillValue = -128b ;
		alloc_greenhouse:long_name = "alloc_greenhouse" ;
		alloc_greenhouse:units = "m3" ;
		alloc_greenhouse:coordinates = "lon lat" ;
		alloc_greenhouse:add_offset = 0.f ;
		alloc_greenhouse:scale_factor = 0.01f ;
	float alloc_wm_dw(time, stations) ;
		alloc_wm_dw:_FillValue = -999.f ;
		alloc_wm_dw:long_name = "alloc_wm_dw" ;
		alloc_wm_dw:units = "m3" ;
		alloc_wm_dw:coordinates = "lon lat" ;
	float demand_agric(time, stations) ;
		demand_agric:_FillValue = -999.f ;
		demand_agric:long_name = "demand_agric" ;
		demand_agric:units = "m3" ;
		demand_agric:coordinates = "lon lat" ;
	float demand_wm(time, stations) ;
		demand_wm:_FillValue = -999.f ;
		demand_wm:long_name = "demand_wm" ;
		demand_wm:units = "m3" ;
		demand_wm:coordinates = "lon lat" ;
	float demand_flush(time, stations) ;
		demand_flush:_FillValue = -999.f ;
		demand_flush:long_name = "demand_flush" ;
		demand_flush:units = "m3" ;
		demand_flush:coordinates = "lon lat" ;
	float demand_flushreturn(time, stations) ;
		demand_flushreturn:_FillValue = -999.f ;
		demand_flushreturn:long_name = "demand_flushreturn" ;
		demand_flushreturn:units = "m3" ;
		demand_flushreturn:coordinates = "lon lat" ;
	byte demand_pubwat(time, stations) ;
		demand_pubwat:_FillValue = -128b ;
		demand_pubwat:long_name = "demand_pubwat" ;
		demand_pubwat:units = "m3" ;
		demand_pubwat:coordinates = "lon lat" ;
		demand_pubwat:add_offset = 0.f ;
		demand_pubwat:scale_factor = 0.01f ;
	byte demand_industry(time, stations) ;
		demand_industry:_FillValue = -128b ;
		demand_industry:long_name = "demand_industry" ;
		demand_industry:units = "m3" ;
		demand_industry:coordinates = "lon lat" ;
		demand_industry:add_offset = 0.f ;
		demand_industry:scale_factor = 0.01f ;
	byte demand_greenhouse(time, stations) ;
		demand_greenhouse:_FillValue = -128b ;
		demand_greenhouse:long_name = "demand_greenhouse" ;
		demand_greenhouse:units = "m3" ;
		demand_greenhouse:coordinates = "lon lat" ;
		demand_greenhouse:add_offset = 0.f ;
		demand_greenhouse:scale_factor = 0.01f ;
	float demand_wmtot(time, stations) ;
		demand_wmtot:_FillValue = -999.f ;
		demand_wmtot:long_name = "demand_wmtot" ;
		demand_wmtot:units = "m3" ;
		demand_wmtot:coordinates = "lon lat" ;
	float demand_wm_todw(time, stations) ;
		demand_wm_todw:_FillValue = -999.f ;
		demand_wm_todw:long_name = "demand_wm_todw" ;
		demand_wm_todw:units = "m3" ;
		demand_wm_todw:coordinates = "lon lat" ;
	float balancecheck(time, stations) ;
		balancecheck:_FillValue = -999.f ;
		balancecheck:long_name = "balancecheck" ;
		balancecheck:units = "m3" ;
		balancecheck:coordinates = "lon lat" ;
// global attributes:
		:Conventions = "CF-1.6" ;
		:title = "LHM parameters van Mozart" ;
		:institution = "Deltares" ;
		:source = "Export archive from Delft-FEWS" ;
		:history = "2018-09-27 06:02:21 GMT: exported from Delft-FEWS" ;
		:references = "http://www.delft-fews.com" ;
		:comment = "Deelgebied=zoetwater; Scenario=Referentie2017" ;
		:Metadata_Conventions = "Unidata Dataset Discovery v1.0" ;
		:summary = "LHM parameters van Mozart" ;
		:date_created = "2018-09-27 06:02:21 GMT" ;
		:Deelgebied = "zoetwater" ;
		:Scenario = "Referentie2017" ;
		:WhatIfScenario = "%WHAT_IF_NAME%" ;
		:fews_implementation_version = "2016.02" ;
		:fews_build_number = "71502" ;
		:fews_patch_number = "68073" ;
		:coordinate_system = "Rijks Driehoekstelsel" ;
		:featureType = "timeSeries" ;
		:time_coverage_start = "1911-01-01T00:00:00+0000" ;
		:time_coverage_end = "1912-01-01T00:00:00+0000" ;
		:geospatial_lon_min = "3.645612377462325" ;
		:geospatial_lon_max = "7.135131693517842" ;
		:geospatial_lat_min = "50.824671652404646" ;
		:geospatial_lat_max = "53.42692119833676" ;
}
